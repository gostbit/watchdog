`ifndef RKV_WATCHDOG_VIRTUAL_SEQUENCER_SV
`define RKV_WATCHDOG_VIRTUAL_SEQUENCER_SV

class rkv_watchdog_virtual_sequencer extends uvm_sequencer;

  rkv_watchdog_config cfg;
  apb_master_sequencer apb_mst_sqr;
  

  `uvm_component_utils(rkv_watchdog_virtual_sequencer)

  function new (string name = "rkv_watchdog_virtual_sequencer", uvm_component parent);
    super.new(name, parent);
  endfunction

  function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    if(!uvm_config_db#(rkv_watchdog_config)::get(this, "", "cfg", cfg)) begin
      `uvm_fatal("GETCFG", "cannot get config object from config DB")
    end
  endfunction



endclass





`endif //RKV_WATCHDOG_VIRTUAL_SEQUENCER_SV
